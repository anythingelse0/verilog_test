module world ();
    wire force = 1'b1;

initial
begin
    $display("Hello,world! %d\n",force);
    
end
endmodule
