module world ();
initial
begin
    $display("Hello,world!");
end
endmodule
